MATLAB 5.0 MAT-file, Platform: PCWIN64, Created on: Wed May 20 09:58:41 2015                                                 IM   U  x��c``������9 4�B�V@�Č@������^�̀D �
�փ�&P�J�A�G(��w��=�|o(�B;@�!� �|T>*���GB���I�A*T>B+�@��Ch�B��"P�W
�ʡ�+!�*�95zC-Լz�y�P��@�k���5�j^Լ�y�P��!t���!�(}`���g
���
�J���w:T_�����f���MS��*��O[r[�;L�N�˞�`|a���i��4�ղ$Mw0h��'9v���]�S������̋���l�T����|�;lC�;D���8ݡ�]���Q��􊧓��8�;  �c 